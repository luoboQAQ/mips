`timescale 1ns/10ps //�� verilog ����û��Ĭ��timescale �ģ�һ��û��ָ�� timescale �� verilog ģ����п��ܴ���ļ̳���ǰ�����ģ�����Чtimescale ������
// �� �� �� �� �� ÿ ��module ��ǰ��ָ��`timescale,timescale �÷���鿴�̲ġ�
`include "ctrl_encode_def.v" //���� C ���Եİ���ͷ�ļ���������Ҳ�����Ƶ�
module mips(clk, reset,out);//�����ļ�
input clk;//�������룬ʱ��Ƶ��
input reset;//�������룬��λ�ź�
output [15:0]out;//�������
assign out=0;
//���������ͱ���
wire [31:2] PC;//��ǰָ���ַ
wire [31:2] NPC;//��һ��ָ���ַ
wire [31:0] Instr;//ָ��
wire [31:0] gpr_read1;//ͨ�üĴ���������RD1 ����
wire [31:0] gpr_read2;//RD2 ����
wire [31:0] Imme32;//�� 16 λ��������չ�õ��� 32 λ������
wire [31:0] ALU_A,A;//ALU ��ԭ������ A
wire [31:0] ALU_B,B;//ALU ��ԭ������ B
wire [31:0] alu_output;//ALU ������
wire [4:0] waddr;//�洢���Ĵ����еĵ�ַ
wire [31:0] inputdata;//�洢������
wire [2:0] NPCOp;//��һ��ָ���ַ�仯���Ϳ����ź�
wire [1:0]EXTOp;//��չ���Ϳ����ź�
wire ASel;//A ������ѡ�����Ϳ����ź�
wire BSel;//B ������ѡ�����Ϳ����ź�
wire [4:0] ALUOp,ALU_ALUOp;
wire Zero;//�ж��Ƿ�Ϊ��ָ֧��
wire [2:0]WDSel;//ͨ�üĴ���д����ѡ������ź�
wire RFWr;//ͨ�üĴ���дʹ�ܿ����ź�
wire [1:0]GPRSel;//ͨ�üĴ���д��ַѡ������ź�
wire [5:0] OP;//opcode
wire [4:0] RS;//ָ�������� rs �ֶ�
wire [4:0] RT;//ָ�������� rt �ֶ�
wire [4:0] RD;//ָ�������� rd �ֶ�
wire [4:0] Shamt;//��λ������ shamt �ֶ�
wire [5:0] Funct;//funct
wire [15:0] Imme16;//16 λ������
wire [25:0] Addr26;//26 λ��ַ
wire nop;
assign OP = Instr[31:26];
assign RS = Instr[25:21];
assign RT = Instr[20:16];
assign RD = Instr[15:11];
assign Shamt = Instr[10:6];
assign Funct = Instr[5:0];
assign Imme16 = Instr[15:0];
assign Addr26 = Instr[25:0];
assign nop =(Instr== 32'b0);
/* main framework of mips-lite-2 *///�����൱�ں�������
pc mips_pc(
       .NPC(NPC),
       .Clk(clk),
       .Reset(reset),
       .PC(PC)
   );//�ṩ pc ��ָ��洢��ȡ��ַ
npc mips_npc(
        .PC(PC),
        .NPCOp(NPCOp),
        .IMM(Addr26),
        .NPC(NPC)
    );//������һ��ָ���ַ�ı仯
im_4k mips_im_4k(
          .addr(PC[11:2]),
          .dout(Instr)
      );//�ṩָ��
ctrl mips_ctrl(
         .opcode(OP),
         .funct(Funct),
         .rt(RT),
         .nop(nop),
         .Zero(Zero),
         .RFWr(RFWr),
         .ALUOp(ALUOp),
         .NPCOp(NPCOp),
         .BSel(BSel),
         .EXTOp(EXTOp),
         .ASel(ASel),
         .GPRSel(GPRSel),
         .WDSel(WDSel)
     );//�������ģ��
gpr mips_gpr(
        .clk(clk),
        .reset(reset),
        .we(RFWr),
        .addr1(RS),
        .addr2(RT),
        .addr3(waddr),
        .inputdata(inputdata),
        .RD1(gpr_read1),
        .RD2(gpr_read2)
    );//ͨ�üĴ���
mux4 MUX_RPR_WD(
         .d0(alu_output),
         .d1(32'b0),
         .d2({PC+1,2'd0}),
         .s(WDSel),
         .y(inputdata)
     );//ѡ������
mux4 MUX_GPR_WA(
         .d0(RD),
         .d1(RT),
         .d2(5'd31),
         .d3(5'd0),
         .s({GPRSel}),
         .y(waddr)
     );//ѡ���ַ
mux2 MUX_ALU_A(
         .d0(gpr_read1),
         .d1({27'd0,Shamt}),
         .s(ASel),
         .y(A)
     );//d1 Ϊ��λ��
mux2 MUX_ALU_B(
         .d0(gpr_read2),
         .d1(Imme32),
         .s(BSel),
         .y(B)
     );
Extend EXTEND(
           .Imm16(Imme16),
           .EXTOp(EXTOp),
           .Imm32(Imme32)
       );//������չ
/*
*ALU ǰ����ʹ ALU ִ����ȷ�Ĳ���
*/
alu_p mips_alu_32_p(
          .A_i(A),
          .B_i(B),
          .ALUOp_i(ALUOp),
          .A_o(ALU_A),
          .B_o(ALU_B),
          .ALUOp_o(ALU_ALUOp)
      );
alu_32 mips_alu_32(
           .A(ALU_A),//.A(A),no
           .B(ALU_B),//.B(B),no
           .ALUOp(ALU_ALUOp),//.ALUOp(ALUOp),no
           .C(alu_output),
           .Zero(Zero)
       );
endmodule