`timescale 1ns/10ps
module gpr(clk, reset, we, addr1, addr2, addr3,inputdata, RD1, RD2);//���� gpr ͨ�üĴ���ģ�飬��ͨ�üĴ����д�ȡ����
input clk;
input reset;//�����ź�
input we;//�ӿ��Ƶ�Ԫ���Ķ�д�����ź�
input [4:0] addr1;//rs
input [4:0] addr2;//rt
input [4:0] addr3;//rd
input [31:0] inputdata;//����[rd]������
output [31:0] RD1;//[rs]����
output [31:0] RD2;//[rt]����
reg [31:0] registers [31:0]; //�Ĵ����ѵ�ʵ��
integer i = 0;
/*
*���� addr3==addr1||addr3==addr2 ʱ�����RD1,RD2 ����
*/
assign RD1 =(clk==1)?registers[addr1]:RD1; //�ӼĴ����ж�Ӧ��ַ addr1 ��λ��ȡ���ݵ� RD1
assign RD2 =(clk==1)?registers[addr2]:RD2; //�ӼĴ����ж�Ӧ��ַ addr2 ��λ��ȡ���ݵ� RD2
/*
��ʼ���Ĵ���
*/
initial begin
    for(i = 0; i < 32; i = i + 1) begin
        registers[i] = 32'h00000000;
    end
end
always @ ( posedge reset or negedge clk) begin//�͵�ƽ��������
    if(reset) begin //����Ƿ�λ�������λ�����³�ʼ���Ĵ����ѣ����򽫽������ addr3��ַ��Ӧ�ļĴ���
        for(i = 0; i <32; i = i + 1) begin
            registers[i] = 32'h00000000;
        end
    end
    else if(we & addr3 != 5'h00) begin //�� 0 �żĴ������ɱ�����
        registers[addr3] <= inputdata;//rd
        // $display("addr: %d, data: %4h",addr3, inputdata);
    end
end
endmodule